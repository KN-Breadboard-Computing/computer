module cpu (
);
    `include "cpu/signals.v"
endmodule
