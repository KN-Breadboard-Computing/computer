module cpu (
    
);
    

endmodule
