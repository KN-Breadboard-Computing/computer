module alu (
    
);
    

endmodule
